module firebird

pub struct Rows {
}
