module firebird

pub struct Result {
pub:
	num_rows_affected int
}
