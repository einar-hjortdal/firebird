module firebirdsql

