module firebird
