module firebird

pub struct Null {}
