module firebird

interface Value {}

// i64
// f64
// bool
// []u8
// string
// time.Time
