module firebird

pub struct Null {}

pub struct NotNull {}
